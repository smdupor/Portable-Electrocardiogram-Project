module heartrate(input clock, input heartbeat, output [7:0] rate);



endmodule